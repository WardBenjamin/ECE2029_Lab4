`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/14/2018 07:26:22 PM
// Design Name: 
// Module Name: mycounter
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mycounter(input clk, output [1:0] Q);
    reg[1:0] temp = 0;
    always @(posedge clk) begin
        temp = temp + 1;
    end
    assign Q = temp;
endmodule
